    Mac OS X            	   2  �     �                                    ATTR;���  �   �                    �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b46827a;Cyberduck;134C74D0-BCDC-4CEC-92C9-2528C14681C1bplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/ipbus-firmware/components/ipbus_slaves/firmware/hdl/ipbus_freq_ctr.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��