    Mac OS X            	   2  �     �                                    ATTR;���  �   �  
                  �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b468277;Cyberduck;605DB49F-7248-4FFD-A46B-2E994D45C307bplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/ipbus-firmware/components/ipbus_core/firmware/hdl/udp_rxram_mux.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             This resource fork intentionally left blank                                                                                                                                                                                                                            ��