    Mac OS X            	   2  �     �                                    ATTR;���  �   �   �                  �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b46825c;Cyberduck;79658ED8-A0A0-4480-87F7-F0F022269828bplist00�_zsftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/neo430/rtl/core/neo430_cfu.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��