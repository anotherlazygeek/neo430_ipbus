    Mac OS X            	   2  �     �                                    ATTR;���  �   �   �                  �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b46825c;Cyberduck;F0900BC2-FA4E-44CA-BEDA-37DF4E195D13bplist00�_zsftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/neo430/rtl/core/neo430_alu.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��