    Mac OS X            	   2  �     �                                    ATTR;���  �   �                    �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b4682a6;Cyberduck;57811F77-25D3-4084-9587-6C286C231D69bplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/ipbus-firmware/boards/glib_v3/base_fw/sim/firmware/hdl/top.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��