    Mac OS X            	   2  �     �                                    ATTR;���  �   �                    �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b468278;Cyberduck;0935CE57-A5BB-4AE5-B2EF-19E51C4210A1bplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/ipbus-firmware/components/ipbus_slaves/firmware/hdl/ipbus_ctr.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               This resource fork intentionally left blank                                                                                                                                                                                                                            ��