    Mac OS X            	   2  �     �                                    ATTR;���  �   �                    �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b468274;Cyberduck;2B253329-D38E-479B-B0BD-490D0F9041EBbplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/ipbus-firmware/components/ipbus_core/firmware/hdl/udp_dualportram_rx.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        This resource fork intentionally left blank                                                                                                                                                                                                                            ��