    Mac OS X            	   2  �     �                                    ATTR;���  �   �  	                  �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b468298;Cyberduck;7918ADF8-8080-4EF0-9AAD-BCC24EFEA141bplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/neo430_ipbus/components/ipbus_core/firmware/hdl/udp_rxram_shim.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              This resource fork intentionally left blank                                                                                                                                                                                                                            ��