    Mac OS X            	   2  �     �                                    ATTR;���  �   �                    �   <  com.apple.quarantine      �  %com.apple.metadata:kMDItemWhereFroms 0081;5b46829d;Cyberduck;65390200-A2F5-401B-9983-9B4645A0CEF6bplist00�_�sftp://excession.phy.bris.ac.uk/usersc/ng18731/ATFC_IPBus_neo_test/neo430_test/myFwArea/src/timing-board-firmware/projects/test/reflect/firmware/hdl/fmc_mirror.vhd
                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         This resource fork intentionally left blank                                                                                                                                                                                                                            ��